module hamming_decoder_precompute(
	input [20:0] ip,
	output reg [15:0] op,
   output reg [4:0] p
	);
reg [20:0] e;
reg a,b,c,d,q,f,g,h,i,j,k,l,m,n,o,r;

always @(ip) begin
e=ip;

a=e[2]^e[6];//
b=e[3]^e[4];//
c=e[7]^e[8];
d=e[15]^e[17]^e[19];
q=e[0]^e[4];//
f=e[1]^e[5];//
g=e[5]^e[6];//
h=e[9]^e[10];
i=e[8]^e[10];//
j=e[9]^e[10];//
k=e[11]^e[12];//
l=e[16]^e[18]^e[20];
m=e[12]^e[14];
n=e[13]^e[14];//
o=e[17]^e[18];//
r=e[19]^e[20];//

p[0]=a^q^i^m^l;
p[1]=a^f^h^n^o;
p[2]=b^g^k^n^r;
p[3]=c^h^k^n;
p[4]=d^l;
case(p) 

5'd3: begin 
op[0]=~e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=e[20];
end
5'd5: begin
op[0]=e[2];
op[1]=~e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=e[20];
end
5'd6: begin
op[0]=e[2];
op[1]=e[4];
op[2]=~e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=e[20];
end

5'd7: begin
	
op[0]=e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=~e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=e[20];
end

5'd9: begin
	
op[0]=e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=~e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=e[20];
end

5'd10: begin
	
op[0]=e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=~e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=e[20];
end

5'd11: begin
	
op[0]=e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=~e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=e[20];
end

5'd12: begin
	
op[0]=e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=~e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=e[20];
end

5'd13: begin
	
op[0]=e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=~e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=e[20];
end

5'd14: begin
	
op[0]=e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=~e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=e[20];
end

5'd15: begin
	
op[0]=e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=~e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=e[20];
end
5'd17: begin
	
op[0]=e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=~e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=e[20];
end

5'd18: begin
	
op[0]=e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=e[16];
op[12]=~e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=e[20];
end

5'd19: begin
	
op[0]=e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=~e[18];
op[14]=e[19];
op[15]=e[20];
end

5'd20: begin
	
op[0]=e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=~e[19];
op[15]=e[20];
end

5'd21: begin
	
op[0]=e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=~e[20];
end

5'd0: begin
op[0]=e[2];
op[1]=e[4];
op[2]=e[5];
op[3]=e[6];
op[4]=e[8];
op[5]=e[9];
op[6]=e[10];
op[7]=e[11];
op[8]=e[12];
op[9]=e[13];
op[10]=e[14];
op[11]=e[16];
op[12]=e[17];
op[13]=e[18];
op[14]=e[19];
op[15]=e[20];
end

endcase
end
endmodule
//010100111100001101100
