module hamming_decoder_serial(
	input [20:0] e,
	input clk,
	output reg [15:0] op,
    output reg [4:0] p
	);
reg [4:0] i;
initial p=0;
initial i=1;
always @ (clk) begin
	if(i==22) begin	
	case(p) 
	
	5'd3: begin 
	op[0]=~e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=e[20];
	end
	5'd5: begin
	op[0]=e[2];
	op[1]=~e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=e[20];
	end
	5'd6: begin
	op[0]=e[2];
	op[1]=e[4];
	op[2]=~e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=e[20];code word 
	end

	5'd7: begin
		
	op[0]=e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=~e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=e[20];
	end

	5'd9: begin
		
	op[0]=e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=~e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=e[20];
	end

	5'd10: begin
		
	op[0]=e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=~e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=e[20];
	end

	5'd11: begin
		
	op[0]=e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=~e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=e[20];
	end

	5'd12: begin
		
	op[0]=e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=~e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=e[20];
	end

	5'd13: begin
		
	op[0]=e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=~e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=e[20];
	end

	5'd14: begin
		
	op[0]=e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=~e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=e[20];
	end

	5'd15: begin
		
	op[0]=e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=~e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=e[20];
	end
	5'd17: begin
		
	op[0]=e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=~e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=e[20];
	end

	5'd18: begin
		
	op[0]=e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=e[16];
	op[12]=~e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=e[20];
	end

	5'd19: begin
		
	op[0]=e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=~e[18];
	op[14]=e[19];
	op[15]=e[20];
	end

	5'd20: begin
		
	op[0]=e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=~e[19];
	op[15]=e[20];
	end

	5'd21: begin	
	op[0]=e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=~e[20];
	end

	5'd0: begin
	op[0]=e[2];
	op[1]=e[4];
	op[2]=e[5];
	op[3]=e[6];
	op[4]=e[8];
	op[5]=e[9];
	op[6]=e[10];
	op[7]=e[11];
	op[8]=e[12];
	op[9]=e[13];
	op[10]=e[14];
	op[11]=e[16];
	op[12]=e[17];
	op[13]=e[18];
	op[14]=e[19];
	op[15]=e[20];
	end

	endcase
	
	end

	else begin
		if(i[0]==1) p[0]=p[0]^e[i-1];
		if(i[1]==1) p[1]=p[1]^e[i-1];
		if(i[2]==1) p[2]=p[2]^e[i-1];
		if(i[3]==1) p[3]=p[3]^e[i-1];
		if(i[4]==1) p[4]=p[4]^e[i-1];
		i=i+1;
	end
end
endmodule
